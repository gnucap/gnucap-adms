
options language=verilog

module foo(1 2);
definedinspice #(.dummy(0)) inst(1 2);
endmodule
